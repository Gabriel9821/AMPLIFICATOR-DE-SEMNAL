** Profile: "SCHEMATIC1-timp"  [ d:\pac\schemaproiect-schematic1-timp.sim ] 

** Creating circuit file "schemaproiect-schematic1-timp.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 1us 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\schemaproiect-SCHEMATIC1.net" 


.END
