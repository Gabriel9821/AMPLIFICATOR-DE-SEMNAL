** Profile: "SCHEMATIC1-frecv"  [ d:\pac\schemaproiect-schematic1-frecv.sim ] 

** Creating circuit file "schemaproiect-schematic1-frecv.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1 500kHz
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\schemaproiect-SCHEMATIC1.net" 


.END
